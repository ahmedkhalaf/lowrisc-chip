// See LICENSE for license details.

module keeper
   (
    input                    clk, rstn,
    nasti_channel            nasti
    );
   
endmodule // keeper
